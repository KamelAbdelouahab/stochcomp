module sadd();

endmodule